*Simulacao

*Alimentacao
Vdd	vdd	0	10
Vss	0	vss	10

*Vin	in	0	AC	1m
*Vin	in	0	SIN(0	1.5	300)
Vin	in	0	1

Rg	in	10	50
R2	10	11	10

Q1	vdd	11	12	Q2N3055
Q2	vss	11	12	QMJ2955

R1	12	0	10

.INCLUDE	2N3055.LIB
.INCLUDE	MJ2955.LIB
.DC	Vin	-10	10	.01

*.TRAN		.1	10	UIC
*.TRAN 1m 2000m 200m 
*.AC	DEC 	1k	.01	1k



.control
run
plot v(12)
set hcopydevtype=postscript
set hcopypscolor=1
hardcopy plot.ps v(12)
.endc


.end
