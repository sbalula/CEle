*Simulacao

*Alimentacao
Vdd	vdd	0	8	
Vss	0	vss	8

*Vin	in	0	AC	1m
*Vin	in	0	SIN(0	1.5	300)
Vin	in	0	1

Rg	in	10	50
R3	10	11	10

Q1	vdd	11	12	Q2N3055
Rsmall	12	121	.001
Q2	121	13	vss	Q2N3055
Q3	13	13	vss	Q2N3055

R2	13	0	10
Rl	12	0	10

.INCLUDE	2N3055.LIB
.DC	Vin	-16	16	.01



*.TRAN		.1	10	UIC
*.TRAN 1m 2000m 200m 
*.AC	DEC 	1k	.01	1k



*.control
*run
*plot v(12), v(out), v(13)
*set hcopydevtype=postscript
*set hcopypscolor=1
*hardcopy plot.ps v(12), v(out), v(13)
*.endc


.end
